`timescale 1ns / 1ps

module FP_MAC_tb();

reg[15:0] A1,A2,A3,A4,A5,A6,A7,A8,A9,A10,A11,A12;
reg [15:0] B1,B2,B3,B4,B5,B6,B7,B8,B9,B10,B11,B12;
reg clk, rst;
wire [15:0] sum;

parameter PERIOD = 1;

FP_MAC test(.rst(rst), .clk(clk),   .A1_x76(A1), .B1_x76(B1), //.P1(P1),
                                    .A2_x76(A2), .B2_x76(B2), //.P2(P2),
                                    .A3_x76(A3), .B3_x76(B3), //.P3(P3),
                                    .A4_x76(A4), .B4_x76(B4), //.P4(P4),
                                    .A5_x76(A5), .B5_x76(B5), //.P5(P5),
                                    .A6_x76(A6), .B6_x76(B6), //.P6(P6),
                                    .A7_x76(A7), .B7_x76(B7), //.P7(P7),
                                    .A8_x76(A8), .B8_x76(B8), //.P8(P8),
                                    .A9_x76(A9), .B9_x76(B9), //.P9(P9),
                                    .A10_x76(A10), .B10_x76(B10), //.P10(P10),
                                    .A11_x76(A11), .B11_x76(B11), //.P11(P11),
                                    .A12_x76(A12), .B12_x76(B12), //.P12(P12)
                                    .sum(sum)
                                    );

initial begin
    clk = 1;
    forever #PERIOD clk = ~clk;
end

initial begin
    rst <= 1; 
    //A <= 16'b0;
    //B <= 16'b0;
    #4;    rst <= 0;
            A1 <= 16'b0_01011_1001100110;    //A = 0.1
            B1 <= 16'b0_01110_0001100110;    //B = 0.55
            
    //#8;    rst <= 1;   #2;     rst <= 0;    
            A2 <= 16'b0_01100_1001100110;    //A = 0.2
            B2 <= 16'b1_01101_1001100110;    //B = -0.4
            
    //#8;    rst <= 1;   #2;     rst <= 0; 
            A3 <= 16'b0_01101_0000000000;    //A = 0.25
            B3 <= 16'b0_01101_0000000000;    //B = 0.25
            
    //#8;    rst <= 1;   #2;     rst <= 0;         
            A4 <= 16'b1_01101_0011001101;    //A = -0.3
            B4 <= 16'b0_01100_0011001101;    //B = 0.15
            
    //#8;     rst <= 1;   #2;     rst <= 0;        
            A5 <= 16'b0_01101_1001100110;    //A = 0.4
            B5 <= 16'b0_01110_0011001101;    //B = 0.6
            
    //#8;      rst <= 1;   #2;     rst <= 0;      
            A6 <= 16'b0_01110_0000000000;    //A = 0.5
            B6 <= 16'b0_01101_1001100110;    //B = 0.4
            
    //#8;     rst <= 1;   #2;     rst <= 0;      
            A7 <= 16'b0_01110_0001100110;    //A = 0.55
            B7 <= 16'b1_01110_1000000000;    //B = -0.75
            
    //#8;     rst <= 1;   #2;     rst <= 0;     
            A8 <= 16'b0_01110_0011001101;    //A = 0.6
            B8 <= 16'b0_01110_1100000000;    //B = 0.875
            
    //#8;     rst <= 1;   #2;     rst <= 0;     
            A9 <= 16'b1_01110_1000000000;    //A = -0.75
            B9 <= 16'b0_01110_1001100110;    //B = 0.8

    //#8;     rst <= 1;   #2;     rst <= 0;     
            A10 <= 16'b0_01110_1001100110;    //A = 0.8
            B10 <= 16'b0_01100_0000000000;    //B = 0.125

    //#8;     rst <= 1;   #2;     rst <= 0;     
            A11 <= 16'b0_01110_1100000000;    //A = 0.875
            B11 <= 16'b1_01110_1110011010;    //B = -0.95

    //#8;     rst <= 1;   #2;     rst <= 0;     
            A12 <= 16'b0_01110_1100110011;    //A = 0.9
            B12 <= 16'b0_01101_0001010010;    //B = 0.27
            
    #100; $finish;
end
endmodule
